module mips_tb();
reg clk1,clk2;
integer k;


mips32 mips32(clk1,clk2);
initial begin
clk1=0; 
clk2=0;
repeat(20)
begin
#5 clk1=1 ;
#5 clk2=0;
#5 clk1=1 ;
#5 clk2=0;
end
end
initial begin
for(k=0;k<31;k=k+1)
mips32.REG[k]=k;

mips32.MEM[0]=32'h2801000a;// addi r1,r0,10
mips32.MEM[1]=32'h28020014;// addi r2,r0,20
mips32.MEM[2]=32'h28030019;// addi r3,r0,30
mips32.MEM[3]=32'h0ce77800;// or r7,r7,r7
mips32.MEM[4]=32'h0ce77800;// or r7,r7,r7
mips32.MEM[5]=32'h00222000;// add r4,r1,r2
mips32.MEM[6]=32'h0ce77800;// or r7,r7,r7
mips32.MEM[7]=32'h00832800;// add r5,r4,r3
mips32.MEM[8]=32'hfc000000;// HLT

mips32.HALTED=0;
mips32.PC=0;
mips32.TAKEN_BRANCH=0;

#280;
for(k=0;k<6;k=k+1)
$display("R%1d - %2d",k,mips32.REG[k]);
#300 $finish;
end
endmodule

module mips32(clk1,clk2);
input clk1,clk2;

reg [31:0] PC,IF_ID_IR,IF_ID_NPC;

reg [31:0] ID_EX_IR,ID_EX_NPC,ID_EX_A,ID_EX_B,ID_EX_Imm;

reg [2:0] ID_EX_TYPE,EX_MEM_TYPE,MEM_WB_TYPE;

reg [31:0] EX_MEM_IR,EX_MEM_ALUOUT,EX_MEM_B;

reg EX_MEM_COND;

reg [31:0] MEM_WB_IR,MEM_WB_ALUOUT,MEM_WB_LMD;

reg [31:0] REG [0:31];

reg [31:0] MEM [0:1023];

parameter ADD=6'b0,SUB=6'b1,AND=6'b10,OR=6'b11,SLT=6'b100,MUL=6'b101,HLT=6'b111111,LW=6'b1000,SW=6'b1001,ADDI=6'b1010,SUBI=6'b1011,SLTI=6'b1100,BNEQZ=6'b1101,BEQZ=6'b1110;

parameter RR_ALU=3'b000,RM_ALU=3'b001,LOAD=3'b010,STORE=3'b011,BRANCH=3'b100,HALT=3'b101;

reg HALTED;
 reg TAKEN_BRANCH;

always @(posedge clk1)// IF STAGE 
if(HALTED==0)
begin
if(((EX_MEM_IR[31:26]==BEQZ) && (EX_MEM_COND ==1)) ||((EX_MEM_IR[31:26]==BNEQZ) && (EX_MEM_COND ==0)))
begin
IF_ID_IR <= #2 MEM[EX_MEM_ALUOUT];
TAKEN_BRANCH <= #2 1'b1;
IF_ID_NPC <= #2 EX_MEM_ALUOUT +1;
PC <= #2 EX_MEM_ALUOUT +1;
end
else
begin
IF_ID_IR <= #2 MEM[PC];
IF_ID_NPC <= #2 PC +1;
PC <= #2 PC +1;
end
end

always @(posedge clk2)
if(HALTED==0)
begin
if(IF_ID_IR[25:21]==5'b00000) ID_EX_A <= 0;
else ID_EX_A <= #2 REG[IF_ID_IR[25:21]];

if(IF_ID_IR[20:16] == 5'b00000) ID_EX_B <= 0;
else ID_EX_B <= #2 REG[IF_ID_IR[20:16]];

ID_EX_NPC <= #2 IF_ID_NPC;
ID_EX_IR <= #2 IF_ID_IR;
ID_EX_Imm <= #2 {{16{IF_ID_IR[15]}},{IF_ID_IR[15:0]}};

case(IF_ID_IR[31:26])
ADD,SUB,AND,OR,SLT,MUL: ID_EX_TYPE <= #2 RR_ALU;
ADDI,SUBI,SLTI        : ID_EX_TYPE <= #2 RM_ALU;
LW                    : ID_EX_TYPE <= #2 LOAD;
SW                    : ID_EX_TYPE <= #2 STORE;
BNEQZ ,BEQZ           : ID_EX_TYPE <= #2 BRANCH;
HLT                   : ID_EX_TYPE <= #2 HALT;
default               : ID_EX_TYPE <= #2 HALT;
endcase
end

always@(posedge clk1)
if(HALTED==0)
begin
EX_MEM_TYPE <= #2 ID_EX_TYPE;
EX_MEM_IR <= #2 ID_EX_IR;
TAKEN_BRANCH <= #2 0;

case(ID_EX_TYPE)
RR_ALU: begin
	case(ID_EX_IR[31:26])
	ADD  : EX_MEM_ALUOUT <= #2 ID_EX_A + ID_EX_B;
	SUB  : EX_MEM_ALUOUT <= #2 ID_EX_A - ID_EX_B;
	AND  : EX_MEM_ALUOUT <= #2 ID_EX_A & ID_EX_B;
	OR   : EX_MEM_ALUOUT <= #2 ID_EX_A | ID_EX_B;
	SLT  : EX_MEM_ALUOUT <= #2 ID_EX_A < ID_EX_B;
	MUL  : EX_MEM_ALUOUT <= #2 ID_EX_A * ID_EX_B;
	default : EX_MEM_ALUOUT <= #2 32'bx;
	endcase
	end

RM_ALU : begin
	case(ID_EX_IR[ 31:26])
	ADDI : EX_MEM_ALUOUT <= #2 ID_EX_A + ID_EX_Imm;
 	SUBI : EX_MEM_ALUOUT <= #2 ID_EX_A - ID_EX_Imm;
	SLTI : EX_MEM_ALUOUT <= #2 ID_EX_A < ID_EX_Imm;
	default :EX_MEM_ALUOUT <= #2 32'hx;
	endcase
	end

LOAD,STORE:
	begin
	EX_MEM_ALUOUT <= #2 ID_EX_A + ID_EX_Imm;
	EX_MEM_B      <= #2 ID_EX_B;
	end
BRANCH   :
	begin
	EX_MEM_ALUOUT <= #2 ID_EX_NPC + ID_EX_Imm;
	EX_MEM_COND   <= #2 (ID_EX_A ==0);
	end
endcase
end
endmodule

























  
